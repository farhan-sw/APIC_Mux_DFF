magic
tech sky130A
timestamp 1744367018
<< nwell >>
rect -105 220 85 560
<< nmos >>
rect 0 0 15 100
<< pmos >>
rect 0 240 15 540
<< ndiff >>
rect -45 85 0 100
rect -45 15 -35 85
rect -15 15 0 85
rect -45 0 0 15
rect 15 85 60 100
rect 15 15 30 85
rect 50 15 60 85
rect 15 0 60 15
<< pdiff >>
rect -45 525 0 540
rect -45 455 -35 525
rect -15 455 0 525
rect -45 425 0 455
rect -45 355 -35 425
rect -15 355 0 425
rect -45 325 0 355
rect -45 255 -35 325
rect -15 255 0 325
rect -45 240 0 255
rect 15 525 60 540
rect 15 455 30 525
rect 50 455 60 525
rect 15 425 60 455
rect 15 355 30 425
rect 50 355 60 425
rect 15 325 60 355
rect 15 255 30 325
rect 50 255 60 325
rect 15 240 60 255
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
<< pdiffc >>
rect -35 455 -15 525
rect -35 355 -15 425
rect -35 255 -15 325
rect 30 455 50 525
rect 30 355 50 425
rect 30 255 50 325
<< psubdiff >>
rect -85 85 -45 100
rect -85 15 -75 85
rect -55 15 -45 85
rect -85 0 -45 15
<< nsubdiff >>
rect -85 525 -45 540
rect -85 455 -75 525
rect -55 455 -45 525
rect -85 425 -45 455
rect -85 355 -75 425
rect -55 355 -45 425
rect -85 325 -45 355
rect -85 255 -75 325
rect -55 255 -45 325
rect -85 240 -45 255
<< psubdiffcont >>
rect -75 15 -55 85
<< nsubdiffcont >>
rect -75 455 -55 525
rect -75 355 -55 425
rect -75 255 -55 325
<< poly >>
rect 0 540 15 555
rect 0 190 15 240
rect -40 180 15 190
rect -40 160 -30 180
rect -10 160 15 180
rect -40 150 15 160
rect 0 100 15 150
rect 0 -15 15 0
<< polycont >>
rect -30 160 -10 180
<< locali >>
rect -35 585 -15 590
rect -35 530 -15 565
rect -85 525 -5 530
rect -85 455 -75 525
rect -55 455 -35 525
rect -15 455 -5 525
rect -85 450 -5 455
rect 20 525 60 530
rect 20 455 30 525
rect 50 455 60 525
rect 20 450 60 455
rect -35 430 -15 450
rect 30 430 50 450
rect -85 425 -5 430
rect -85 355 -75 425
rect -55 355 -35 425
rect -15 355 -5 425
rect -85 350 -5 355
rect 20 425 60 430
rect 20 355 30 425
rect 50 355 60 425
rect 20 350 60 355
rect -35 330 -15 350
rect 30 330 50 350
rect -85 325 -5 330
rect -85 255 -75 325
rect -55 255 -35 325
rect -15 255 -5 325
rect -85 250 -5 255
rect 20 325 60 330
rect 20 255 30 325
rect 50 255 60 325
rect 20 250 60 255
rect 30 190 50 250
rect -40 180 0 190
rect -40 160 -30 180
rect -10 160 0 180
rect -40 150 0 160
rect 30 180 70 190
rect 30 160 40 180
rect 60 160 70 180
rect 30 150 70 160
rect 30 90 50 150
rect -85 85 -5 90
rect -85 15 -75 85
rect -55 15 -35 85
rect -15 15 -5 85
rect -85 10 -5 15
rect 20 85 60 90
rect 20 15 30 85
rect 50 15 60 85
rect 20 10 60 15
rect -35 -25 -15 10
<< viali >>
rect -35 565 -15 585
rect -30 160 -10 180
rect 40 160 60 180
rect -35 -45 -15 -25
<< metal1 >>
rect -105 585 85 590
rect -105 565 -35 585
rect -15 565 85 585
rect -105 560 85 565
rect -40 180 0 190
rect -40 160 -30 180
rect -10 160 0 180
rect -40 150 0 160
rect 30 180 70 190
rect 30 160 40 180
rect 60 160 70 180
rect 30 150 70 160
rect -105 -25 85 -20
rect -105 -45 -35 -25
rect -15 -45 85 -25
rect -105 -50 85 -45
<< labels >>
flabel metal1 -40 150 -40 190 1 FreeSans 200 0 0 0 A
port 1 n
flabel metal1 70 150 70 190 1 FreeSans 200 0 0 0 OUT
port 2 n
flabel metal1 -105 560 -105 590 3 FreeSans 200 0 0 0 VP
port 3 e
flabel metal1 -105 -50 -105 -20 3 FreeSans 200 0 0 0 VN
port 4 e
<< end >>
