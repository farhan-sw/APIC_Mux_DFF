* NGSPICE file created from nand.ext - technology: sky130A

.subckt nand A B OUT VP VN
X0 OUT B a_30_0# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
**devattr s=10000,300 d=20000,600
X1 a_30_0# A VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
**devattr s=18000,580 d=10000,300
X2 OUT A VP VP sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.425 ps=6.95 w=3 l=0.15
**devattr s=54000,1380 d=30000,700
X3 VP B OUT VP sky130_fd_pr__pfet_01v8 ad=1.425 pd=6.95 as=0.75 ps=3.5 w=3 l=0.15
**devattr s=30000,700 d=60000,1400
.ends

