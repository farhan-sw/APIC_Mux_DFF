magic
tech sky130A
magscale 1 2
timestamp 1744416606
<< nwell >>
rect 1270 540 1310 1220
rect 2200 540 2250 1220
<< metal1 >>
rect 0 1220 30 1280
rect 1270 1220 1310 1280
rect 2200 1220 2240 1280
rect 1160 650 1240 660
rect 1160 590 1170 650
rect 1230 640 1240 650
rect 2530 650 2610 660
rect 2530 640 2540 650
rect 1230 600 2540 640
rect 1230 590 1240 600
rect 1160 580 1240 590
rect 2530 590 2540 600
rect 2600 590 2610 650
rect 2530 580 2610 590
rect 510 490 590 530
rect 130 470 210 480
rect 130 460 140 470
rect 40 420 140 460
rect 130 410 140 420
rect 200 410 210 470
rect 130 400 210 410
rect 270 450 590 490
rect 1440 520 1520 530
rect 1160 470 1240 480
rect 270 400 350 450
rect 1160 410 1170 470
rect 1230 410 1240 470
rect 1440 460 1450 520
rect 1510 460 1520 520
rect 2370 490 2450 530
rect 1440 450 1520 460
rect 2090 450 2450 490
rect 2530 520 2610 530
rect 2530 460 2540 520
rect 2600 460 2610 520
rect 2530 450 2610 460
rect 1160 400 1240 410
rect 2090 400 2170 450
rect 3020 400 3100 480
rect 670 360 750 400
rect 40 320 750 360
rect 1600 390 1680 400
rect 1600 330 1610 390
rect 1670 330 1680 390
rect 1600 320 1680 330
rect 1440 310 1520 320
rect 1440 280 1450 310
rect 40 250 1450 280
rect 1510 250 1520 310
rect 40 240 1520 250
rect 1600 190 1680 200
rect 130 170 210 180
rect 130 110 140 170
rect 200 160 210 170
rect 1600 160 1610 190
rect 200 130 1610 160
rect 1670 130 1680 190
rect 200 120 1680 130
rect 200 110 210 120
rect 130 100 210 110
rect 0 0 30 60
rect 1270 0 1310 60
rect 2200 0 2240 60
<< via1 >>
rect 1170 590 1230 650
rect 2540 590 2600 650
rect 140 410 200 470
rect 1170 410 1230 470
rect 1450 460 1510 520
rect 2540 460 2600 520
rect 1610 330 1670 390
rect 1450 250 1510 310
rect 140 110 200 170
rect 1610 130 1670 190
<< metal2 >>
rect 1160 650 1240 660
rect 1160 590 1170 650
rect 1230 590 1240 650
rect 1160 580 1240 590
rect 2530 650 2610 660
rect 2530 590 2540 650
rect 2600 590 2610 650
rect 2530 580 2610 590
rect 1180 480 1220 580
rect 2550 530 2590 580
rect 1440 520 1520 530
rect 130 470 210 480
rect 130 410 140 470
rect 200 410 210 470
rect 130 400 210 410
rect 1160 470 1240 480
rect 1160 410 1170 470
rect 1230 410 1240 470
rect 1440 460 1450 520
rect 1510 460 1520 520
rect 1440 450 1520 460
rect 2530 520 2610 530
rect 2530 460 2540 520
rect 2600 460 2610 520
rect 2530 450 2610 460
rect 1160 400 1240 410
rect 150 180 190 400
rect 1460 320 1500 450
rect 1600 390 1680 400
rect 1600 330 1610 390
rect 1670 330 1680 390
rect 1600 320 1680 330
rect 1440 310 1520 320
rect 1440 250 1450 310
rect 1510 250 1520 310
rect 1440 240 1520 250
rect 1620 200 1660 320
rect 1600 190 1680 200
rect 130 170 210 180
rect 130 110 140 170
rect 200 110 210 170
rect 1600 130 1610 190
rect 1670 130 1680 190
rect 1600 120 1680 130
rect 130 100 210 110
use and  and_0
timestamp 1744378255
transform 1 0 380 0 1 0
box 0 0 931 1280
use and  and_1
timestamp 1744378255
transform 1 0 1310 0 1 0
box 0 0 931 1280
use inverter  inverter_0
timestamp 1744367018
transform 1 0 210 0 1 100
box -210 -100 170 1180
use or  or_0
timestamp 1744376768
transform 1 0 2240 0 1 0
box 0 0 931 1280
<< labels >>
flabel metal1 40 420 40 460 1 FreeSans 400 0 0 0 S
port 3 n
flabel metal1 40 320 40 360 1 FreeSans 400 0 0 0 A
port 1 n
flabel metal1 40 240 40 280 1 FreeSans 400 0 0 0 B
port 2 n
flabel metal1 3100 400 3100 480 1 FreeSans 400 0 0 0 D
port 4 n
flabel metal1 0 1220 0 1280 3 FreeSans 400 0 0 0 VP
port 5 e
flabel metal1 0 0 0 60 3 FreeSans 400 0 0 0 VN
port 6 e
<< end >>
