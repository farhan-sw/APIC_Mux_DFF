** sch_path: /foss/designs/APIC_Mux_DFF/basic_cell/single_cell/inverter/tb_xschem_inverter.sch
**.subckt tb_xschem_inverter A OUT A
*.ipin A
*.opin OUT
*.ipin A
x2 VDD A OUT GND inverter
V3 VDD GND 1.8
V4 A GND pulse(0 1.8 0ns 0.1ns 0.1ns 20ns 40ns)
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt


.control
save all
tran 0.1ns 80ns
plot v(A) v(OUT)+2
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/APIC_Mux_DFF/basic_cell/single_cell/inverter/inverter.sym # of pins=4
** sym_path: /foss/designs/APIC_Mux_DFF/basic_cell/single_cell/inverter/inverter.sym
** sch_path: /foss/designs/APIC_Mux_DFF/basic_cell/single_cell/inverter/inverter.sch
.subckt inverter VP A OUT VN
*.ipin A
*.ipin VP
*.ipin VN
*.opin OUT
XM1 OUT A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
