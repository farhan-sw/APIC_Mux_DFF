* PEX produced on Sat Apr 12 05:42:19 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from mux.ext - technology: sky130A

.subckt mux A B S D VP VN
X0 or_0.nor_0.OUT.t1 or_0.B.t2 a_2480_580.t1 VP.t14 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X1 a_2480_580.t0 or_0.A.t2 VP.t9 VP.t8 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X2 VP.t3 A.t0 and_0.nand_0.OUT.t2 VP.t2 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X3 D.t1 or_0.nor_0.OUT.t3 VN.t17 VN.t16 sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X4 D.t0 or_0.nor_0.OUT.t4 VP.t16 VP.t15 sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X5 or_0.B.t0 and_0.nand_0.OUT.t3 VN.t1 VN.t0 sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X6 or_0.B.t1 and_0.nand_0.OUT.t4 VP.t18 VP.t17 sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X7 and_1.nand_0.OUT.t0 S.t0 a_1550_100.t0 VN.t15 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X8 a_1550_100.t1 B.t0 VN.t9 VN.t8 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X9 or_0.A.t1 and_1.nand_0.OUT.t3 VN.t5 VN.t4 sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X10 VP.t13 S.t1 and_1.nand_0.OUT.t1 VP.t12 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X11 inverter_0.OUT.t1 S.t2 VN.t11 VN.t10 sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X12 and_1.nand_0.OUT.t2 B.t1 VP.t5 VP.t4 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X13 or_0.A.t0 and_1.nand_0.OUT.t4 VP.t1 VP.t0 sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X14 a_620_100.t0 inverter_0.OUT.t2 VN.t3 VN.t2 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X15 inverter_0.OUT.t0 S.t3 VP.t11 VP.t10 sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X16 VN.t14 or_0.B.t3 or_0.nor_0.OUT.t0 VN.t13 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X17 and_0.nand_0.OUT.t0 inverter_0.OUT.t3 VP.t7 VP.t6 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X18 and_0.nand_0.OUT.t1 A.t1 a_620_100.t1 VN.t12 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X19 or_0.nor_0.OUT.t2 or_0.A.t3 VN.t7 VN.t6 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
R0 or_0.B.n0 or_0.B.t2 586.433
R1 or_0.B.n0 or_0.B.t3 425.767
R2 or_0.B.n1 or_0.B.t1 190.534
R3 or_0.B.n1 or_0.B.t0 180.101
R4 or_0.nor_0.B or_0.B.n0 161.3
R5 or_0.nor_0.B or_0.B.n1 32.1755
R6 a_2480_580.t0 a_2480_580.t1 32.8338
R7 or_0.nor_0.OUT.n0 or_0.nor_0.OUT.t4 660.194
R8 or_0.nor_0.OUT.n0 or_0.nor_0.OUT.t3 338.861
R9 or_0.nor_0.OUT.n2 or_0.nor_0.OUT.t1 209.733
R10 or_0.nor_0.OUT or_0.nor_0.OUT.n0 161.363
R11 or_0.nor_0.OUT.n2 or_0.nor_0.OUT.n1 156.5
R12 or_0.nor_0.OUT.n1 or_0.nor_0.OUT.t0 30.0005
R13 or_0.nor_0.OUT.n1 or_0.nor_0.OUT.t2 30.0005
R14 or_0.nor_0.OUT or_0.nor_0.OUT.n2 9.363
R15 VP.t0 VP.n20 384.192
R16 VP.n61 VP.t17 384.192
R17 VP.t14 VP.n11 328.31
R18 VP.n66 VP.t12 328.31
R19 VP.n50 VP.t2 328.31
R20 VP.n45 VP.t10 328.31
R21 VP.n33 VP.n31 300
R22 VP.n27 VP.n26 300
R23 VP.n49 VP.n25 300
R24 VP.n22 VP.n21 300
R25 VP.n65 VP.n2 300
R26 VP.n13 VP.n12 300
R27 VP.n10 VP.n4 300
R28 VP.n36 VP.n35 292.5
R29 VP.n41 VP.n40 292.5
R30 VP.n48 VP.n46 292.5
R31 VP.n57 VP.n56 292.5
R32 VP.n64 VP.n62 292.5
R33 VP.n16 VP.n15 292.5
R34 VP.n9 VP.n5 292.5
R35 VP.n11 VP.t15 202.575
R36 VP.n20 VP.t8 202.575
R37 VP.n66 VP.t0 202.575
R38 VP.t4 VP.n61 202.575
R39 VP.n50 VP.t17 202.575
R40 VP.t6 VP.n45 202.575
R41 VP.n32 VP.t10 202.575
R42 VP.n28 VP.t3 183.833
R43 VP.n23 VP.t13 183.833
R44 VP.t8 VP.t14 181.619
R45 VP.t12 VP.t4 181.619
R46 VP.t2 VP.t6 181.619
R47 VP.n44 VP.n43 149.718
R48 VP.n52 VP.n51 149.718
R49 VP.n60 VP.n59 149.718
R50 VP.n68 VP.n67 149.718
R51 VP.n19 VP.n18 149.718
R52 VP.n36 VP.n29 149.718
R53 VP.n6 VP.n3 149.718
R54 VP.n35 VP.n34 141.603
R55 VP.n42 VP.n41 140.119
R56 VP.n46 VP.n24 140.119
R57 VP.n58 VP.n57 140.119
R58 VP.n62 VP.n1 140.119
R59 VP.n17 VP.n16 140.119
R60 VP.n7 VP.n5 140.119
R61 VP.n34 VP.n33 108.195
R62 VP.n40 VP.n26 98.9005
R63 VP.n49 VP.n48 98.9005
R64 VP.n56 VP.n21 98.9005
R65 VP.n65 VP.n64 98.9005
R66 VP.n15 VP.n12 98.9005
R67 VP.n10 VP.n9 98.9005
R68 VP.n14 VP.n13 92.5005
R69 VP.n20 VP.n12 92.5005
R70 VP.n63 VP.n2 92.5005
R71 VP.n66 VP.n65 92.5005
R72 VP.n55 VP.n22 92.5005
R73 VP.n61 VP.n21 92.5005
R74 VP.n47 VP.n25 92.5005
R75 VP.n50 VP.n49 92.5005
R76 VP.n39 VP.n27 92.5005
R77 VP.n45 VP.n26 92.5005
R78 VP.n31 VP.n30 92.5005
R79 VP.n33 VP.n32 92.5005
R80 VP.n11 VP.n10 92.5005
R81 VP.n8 VP.n4 92.5005
R82 VP.n31 VP.n29 57.2175
R83 VP.n19 VP.n13 57.2175
R84 VP.n67 VP.n2 57.2175
R85 VP.n60 VP.n22 57.2175
R86 VP.n51 VP.n25 57.2175
R87 VP.n44 VP.n27 57.2175
R88 VP.n4 VP.n3 57.2175
R89 VP.n6 VP 44.8338
R90 VP.n37 VP.n36 44.5005
R91 VP.n43 VP.n38 44.5005
R92 VP.n53 VP.n52 44.5005
R93 VP.n59 VP.n54 44.5005
R94 VP.n69 VP.n68 44.5005
R95 VP.n18 VP.n0 44.5005
R96 VP.n36 VP.n30 25.6005
R97 VP.n40 VP.n39 19.2005
R98 VP.n48 VP.n47 19.2005
R99 VP.n56 VP.n55 19.2005
R100 VP.n64 VP.n63 19.2005
R101 VP.n15 VP.n14 19.2005
R102 VP.n9 VP.n8 19.2005
R103 VP.n20 VP.n19 17.6428
R104 VP.n67 VP.n66 17.6428
R105 VP.n61 VP.n60 17.6428
R106 VP.n51 VP.n50 17.6428
R107 VP.n45 VP.n44 17.6428
R108 VP.n32 VP.n29 17.6428
R109 VP.n11 VP.n3 17.6428
R110 VP.n35 VP.t11 16.4172
R111 VP.n41 VP.t7 16.4172
R112 VP.n46 VP.t18 16.4172
R113 VP.n57 VP.t5 16.4172
R114 VP.n62 VP.t1 16.4172
R115 VP.n16 VP.t9 16.4172
R116 VP.n5 VP.t16 16.4172
R117 VP.n43 VP.n42 12.2643
R118 VP.n42 VP.n39 12.2643
R119 VP.n52 VP.n24 12.2643
R120 VP.n47 VP.n24 12.2643
R121 VP.n59 VP.n58 12.2643
R122 VP.n58 VP.n55 12.2643
R123 VP.n68 VP.n1 12.2643
R124 VP.n63 VP.n1 12.2643
R125 VP.n18 VP.n17 12.2643
R126 VP.n17 VP.n14 12.2643
R127 VP.n7 VP.n6 12.2643
R128 VP.n8 VP.n7 12.2643
R129 VP.n34 VP.n30 9.29594
R130 VP VP.n0 0.729667
R131 VP VP.n69 0.542167
R132 VP.n54 VP.n23 0.542167
R133 VP VP.n53 0.542167
R134 VP.n38 VP.n28 0.542167
R135 VP VP.n37 0.458833
R136 VP VP.n0 0.333833
R137 VP.n69 VP 0.333833
R138 VP.n54 VP 0.333833
R139 VP.n53 VP 0.333833
R140 VP.n38 VP 0.333833
R141 VP.n37 VP 0.333833
R142 VP.n23 VP 0.188
R143 VP.n28 VP 0.188
R144 or_0.A.n0 or_0.A.t2 579.861
R145 or_0.A.n0 or_0.A.t3 419.195
R146 or_0.A.n1 or_0.A.t0 190.534
R147 or_0.A.n1 or_0.A.t1 180.101
R148 or_0.nor_0.A or_0.A.n0 161.363
R149 and_1.inverter_0.OUT or_0.A.n1 9.35606
R150 and_1.inverter_0.OUT or_0.nor_0.A 0.6255
R151 A.n0 A.t0 795.301
R152 A.n0 A.t1 216.9
R153 A A.n0 161.363
R154 and_0.nand_0.OUT.n0 and_0.nand_0.OUT.t4 660.194
R155 and_0.nand_0.OUT.n0 and_0.nand_0.OUT.t3 338.861
R156 and_0.nand_0.OUT.n2 and_0.nand_0.OUT.t1 196.101
R157 and_0.nand_0.OUT.n2 and_0.nand_0.OUT.n1 183.718
R158 and_0.nand_0.OUT and_0.nand_0.OUT.n0 161.3
R159 and_0.nand_0.OUT.n1 and_0.nand_0.OUT.t2 16.4172
R160 and_0.nand_0.OUT.n1 and_0.nand_0.OUT.t0 16.4172
R161 and_0.nand_0.OUT and_0.nand_0.OUT.n2 9.363
R162 VN.t4 VN.n5 2240.74
R163 VN.n16 VN.t0 2240.74
R164 VN.t13 VN.n3 1914.81
R165 VN.n17 VN.t15 1914.81
R166 VN.n11 VN.t12 1914.81
R167 VN.n10 VN.t10 1914.81
R168 VN.n6 VN.t10 1772.88
R169 VN.n3 VN.t16 1181.48
R170 VN.n5 VN.t6 1181.48
R171 VN.n17 VN.t4 1181.48
R172 VN.t8 VN.n16 1181.48
R173 VN.n11 VN.t0 1181.48
R174 VN.t2 VN.n10 1181.48
R175 VN.t6 VN.t13 1059.26
R176 VN.t15 VN.t8 1059.26
R177 VN.t12 VN.t2 1059.26
R178 VN.n10 VN.n9 591.4
R179 VN.n12 VN.n11 591.4
R180 VN.n16 VN.n15 591.4
R181 VN.n18 VN.n17 591.4
R182 VN.n5 VN.n4 591.4
R183 VN.n3 VN.n2 591.4
R184 VN.n1 VN.t14 173.4
R185 VN.n6 VN.t11 122.501
R186 VN.n9 VN.t3 122.501
R187 VN.n12 VN.t1 122.501
R188 VN.n15 VN.t9 122.501
R189 VN.n18 VN.t5 122.501
R190 VN.n4 VN.t7 122.501
R191 VN.n2 VN.t17 122.501
R192 VN.n2 VN 38.4338
R193 VN.n7 VN.n6 38.1005
R194 VN.n9 VN.n8 38.1005
R195 VN.n13 VN.n12 38.1005
R196 VN.n15 VN.n14 38.1005
R197 VN.n19 VN.n18 38.1005
R198 VN.n4 VN.n0 38.1005
R199 VN.n14 VN 0.729667
R200 VN.n8 VN 0.729667
R201 VN.n1 VN.n0 0.542167
R202 VN VN.n19 0.542167
R203 VN VN.n13 0.542167
R204 VN VN.n7 0.458833
R205 VN VN.n0 0.333833
R206 VN.n19 VN 0.333833
R207 VN.n14 VN 0.333833
R208 VN.n13 VN 0.333833
R209 VN.n8 VN 0.333833
R210 VN.n7 VN 0.333833
R211 VN VN.n1 0.188
R212 D.n0 D.t0 190.534
R213 D.n0 D.t1 180.101
R214 D D.n0 9.363
R215 S.n0 S.t1 795.301
R216 S.n2 S.t3 660.194
R217 S.n2 S.t2 338.861
R218 S.n0 S.t0 216.9
R219 S.n3 S.n2 161.3
R220 S.n1 S.n0 161.3
R221 S.n3 S.n1 23.7817
R222 S.n1 S 0.063
R223 S S.n3 0.063
R224 a_1550_100.t0 a_1550_100.t1 60.0005
R225 and_1.nand_0.OUT.n0 and_1.nand_0.OUT.t4 660.194
R226 and_1.nand_0.OUT.n0 and_1.nand_0.OUT.t3 338.861
R227 and_1.nand_0.OUT.n2 and_1.nand_0.OUT.t0 196.101
R228 and_1.nand_0.OUT.n2 and_1.nand_0.OUT.n1 183.718
R229 and_1.nand_0.OUT and_1.nand_0.OUT.n0 161.3
R230 and_1.nand_0.OUT.n1 and_1.nand_0.OUT.t1 16.4172
R231 and_1.nand_0.OUT.n1 and_1.nand_0.OUT.t2 16.4172
R232 and_1.nand_0.OUT and_1.nand_0.OUT.n2 9.363
R233 B.n0 B.t1 579.861
R234 B.n0 B.t0 419.195
R235 B.n1 B.n0 161.3
R236 B.n1 B 13.9693
R237 B B.n1 0.063
R238 inverter_0.OUT.n0 inverter_0.OUT.t3 579.861
R239 inverter_0.OUT.n0 inverter_0.OUT.t2 419.195
R240 inverter_0.OUT.n1 inverter_0.OUT.t0 190.534
R241 inverter_0.OUT.n1 inverter_0.OUT.t1 180.101
R242 inverter_0.OUT inverter_0.OUT.n0 161.363
R243 inverter_0.OUT inverter_0.OUT.n1 9.35606
R244 a_620_100.t0 a_620_100.t1 60.0005
C0 S inverter_0.OUT 0.17868f
C1 VP inverter_0.OUT 0.53047f
C2 S and_0.nand_0.OUT 0.03678f
C3 S and_1.nand_0.OUT 0.17419f
C4 and_0.nand_0.OUT VP 0.60492f
C5 and_1.nand_0.OUT VP 0.54461f
C6 D VP 0.23886f
C7 or_0.nor_0.OUT D 0.12966f
C8 and_0.nand_0.OUT inverter_0.OUT 0.08389f
C9 A B 0.35309f
C10 S B 0.66501f
C11 B VP 0.1302f
C12 A S 0.13507f
C13 A VP 0.08326f
C14 B inverter_0.OUT 0.03505f
C15 A inverter_0.OUT 0.23255f
C16 and_0.nand_0.OUT B 0.13927f
C17 S VP 0.21218f
C18 and_1.nand_0.OUT B 0.08079f
C19 A and_0.nand_0.OUT 0.1476f
C20 or_0.nor_0.OUT VP 0.32179f
C21 D VN 0.36092f
C22 B VN 0.6162f
C23 A VN 0.29263f
C24 S VN 1.69147f
C25 VP VN 7.0416f
C26 or_0.nor_0.OUT VN 0.70285f
C27 and_1.nand_0.OUT VN 0.53204f
C28 and_0.nand_0.OUT VN 0.46924f
C29 inverter_0.OUT VN 0.49836f
.ends

