magic
tech sky130A
timestamp 1744388325
<< poly >>
rect 1055 225 1060 265
<< locali >>
rect 1055 225 1060 265
rect 1180 225 1185 265
<< metal1 >>
rect 0 610 15 640
rect 65 325 105 330
rect 65 295 70 325
rect 100 320 105 325
rect 510 325 550 330
rect 510 320 515 325
rect 100 300 515 320
rect 100 295 105 300
rect 65 290 105 295
rect 510 295 515 300
rect 545 295 550 325
rect 510 290 550 295
rect 255 245 295 265
rect 65 235 105 240
rect 65 230 70 235
rect 0 210 70 230
rect 65 205 70 210
rect 100 205 105 235
rect 65 200 105 205
rect 135 225 295 245
rect 380 260 420 265
rect 380 230 385 260
rect 415 230 420 260
rect 380 225 420 230
rect 510 260 550 265
rect 510 230 515 260
rect 545 230 550 260
rect 510 225 550 230
rect 635 245 805 265
rect 635 225 675 245
rect 765 225 805 245
rect 890 245 1060 265
rect 890 225 930 245
rect 1020 225 1060 245
rect 1145 260 1185 265
rect 1145 230 1150 260
rect 1180 230 1185 260
rect 1145 225 1185 230
rect 135 200 175 225
rect 335 180 375 200
rect 845 195 885 200
rect 0 160 590 180
rect 845 165 850 195
rect 880 165 885 195
rect 845 160 885 165
rect 1100 195 1140 200
rect 1100 165 1105 195
rect 1135 165 1140 195
rect 1100 160 1140 165
rect 385 135 425 140
rect 385 105 390 135
rect 420 130 425 135
rect 1100 135 1140 140
rect 1100 130 1105 135
rect 420 110 1105 130
rect 420 105 425 110
rect 385 100 425 105
rect 1100 105 1105 110
rect 1135 105 1140 135
rect 1100 100 1140 105
rect 845 85 885 90
rect 845 55 850 85
rect 880 80 885 85
rect 1165 85 1205 90
rect 1165 80 1170 85
rect 880 60 1170 80
rect 880 55 885 60
rect 845 50 885 55
rect 1165 55 1170 60
rect 1200 55 1205 85
rect 1165 50 1205 55
rect 0 0 15 30
<< via1 >>
rect 70 295 100 325
rect 515 295 545 325
rect 70 205 100 235
rect 385 230 415 260
rect 515 230 545 260
rect 1150 230 1180 260
rect 850 165 880 195
rect 1105 165 1135 195
rect 390 105 420 135
rect 1105 105 1135 135
rect 850 55 880 85
rect 1170 55 1200 85
<< metal2 >>
rect 65 325 105 330
rect 65 295 70 325
rect 100 295 105 325
rect 65 290 105 295
rect 510 325 550 330
rect 510 295 515 325
rect 545 295 550 325
rect 510 290 550 295
rect 75 240 95 290
rect 520 265 540 290
rect 380 260 420 265
rect 65 235 105 240
rect 65 205 70 235
rect 100 205 105 235
rect 380 230 385 260
rect 415 230 420 260
rect 380 225 420 230
rect 510 260 550 265
rect 510 230 515 260
rect 545 230 550 260
rect 510 225 550 230
rect 1145 260 1185 265
rect 1145 230 1150 260
rect 1180 230 1185 260
rect 1145 225 1185 230
rect 65 200 105 205
rect 400 140 420 225
rect 845 195 885 200
rect 845 165 850 195
rect 880 165 885 195
rect 845 160 885 165
rect 1100 195 1140 200
rect 1100 165 1105 195
rect 1135 165 1140 195
rect 1100 160 1140 165
rect 385 135 425 140
rect 385 105 390 135
rect 420 105 425 135
rect 385 100 425 105
rect 855 90 875 160
rect 1110 140 1130 160
rect 1100 135 1140 140
rect 1100 105 1105 135
rect 1135 105 1140 135
rect 1100 100 1140 105
rect 1170 90 1185 225
rect 845 85 885 90
rect 845 55 850 85
rect 880 55 885 85
rect 845 50 885 55
rect 1165 85 1205 90
rect 1165 55 1170 85
rect 1200 55 1205 85
rect 1165 50 1205 55
use inverter  inverter_1
timestamp 1744367018
transform 1 0 105 0 1 50
box -105 -50 85 590
use nand  nand_0
timestamp 1744370894
transform 1 0 295 0 1 50
box -105 -50 150 590
use nand  nand_1
timestamp 1744370894
transform 1 0 550 0 1 50
box -105 -50 150 590
use nand  nand_2
timestamp 1744370894
transform 1 0 1060 0 1 50
box -105 -50 150 590
use nand  nand_3
timestamp 1744370894
transform 1 0 805 0 1 50
box -105 -50 150 590
<< labels >>
flabel metal1 0 210 0 230 3 FreeSans 200 0 0 0 D
port 1 e
flabel metal1 0 160 0 180 3 FreeSans 200 0 0 0 Clk
port 2 e
flabel metal1 0 610 0 640 3 FreeSans 200 0 0 0 VP
port 5 e
flabel metal1 0 0 0 30 3 FreeSans 200 0 0 0 VN
port 6 e
flabel metal1 1060 225 1060 265 1 FreeSans 200 0 0 0 Q
port 3 n
flabel metal2 1185 225 1185 265 1 FreeSans 200 0 0 0 Qi
port 4 n
<< end >>
