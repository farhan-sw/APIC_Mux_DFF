* PEX produced on Sat Apr 12 05:27:26 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from and.ext - technology: sky130A

.subckt and A B OUT VP VN
X0 OUT.t0 nand_0.OUT.t3 VP.t1 VP.t0 sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X1 nand_0.OUT.t2 B.t0 a_240_100.t1 VN.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X2 a_240_100.t0 A.t0 VN.t3 VN.t2 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X3 VP.t3 B.t1 nand_0.OUT.t0 VP.t2 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X4 nand_0.OUT.t1 A.t1 VP.t5 VP.t4 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X5 OUT.t1 nand_0.OUT.t4 VN.t1 VN.t0 sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
R0 nand_0.OUT.n0 nand_0.OUT.t3 660.194
R1 nand_0.OUT.n0 nand_0.OUT.t4 338.861
R2 nand_0.OUT.n2 nand_0.OUT.t2 196.101
R3 nand_0.OUT.n2 nand_0.OUT.n1 183.718
R4 nand_0.OUT nand_0.OUT.n0 161.3
R5 nand_0.OUT.n1 nand_0.OUT.t0 16.4172
R6 nand_0.OUT.n1 nand_0.OUT.t1 16.4172
R7 nand_0.OUT nand_0.OUT.n2 9.363
R8 VP.t2 VP.n11 328.31
R9 VP.n13 VP.n3 300
R10 VP.n10 VP.n5 300
R11 VP.n16 VP.n15 292.5
R12 VP.n9 VP.n6 292.5
R13 VP.n11 VP.t0 202.575
R14 VP.n12 VP.t4 202.575
R15 VP.n18 VP.t3 183.833
R16 VP.t4 VP.t2 181.619
R17 VP.n16 VP.n1 149.718
R18 VP.n4 VP.n0 149.718
R19 VP.n15 VP.n14 141.603
R20 VP.n7 VP.n6 140.119
R21 VP.n14 VP.n13 108.195
R22 VP.n10 VP.n9 98.9005
R23 VP.n3 VP.n2 92.5005
R24 VP.n13 VP.n12 92.5005
R25 VP.n11 VP.n10 92.5005
R26 VP.n8 VP.n5 92.5005
R27 VP.n3 VP.n1 57.2175
R28 VP.n5 VP.n4 57.2175
R29 VP VP.n0 44.8338
R30 VP.n17 VP.n16 44.5005
R31 VP.n16 VP.n2 25.6005
R32 VP.n9 VP.n8 19.2005
R33 VP.n12 VP.n1 17.6428
R34 VP.n11 VP.n4 17.6428
R35 VP.n15 VP.t5 16.4172
R36 VP.n6 VP.t1 16.4172
R37 VP.n7 VP.n0 12.2643
R38 VP.n8 VP.n7 12.2643
R39 VP.n14 VP.n2 9.29594
R40 VP.n18 VP.n17 0.542167
R41 VP.n17 VP 0.333833
R42 VP VP.n18 0.188
R43 OUT.n0 OUT.t0 190.534
R44 OUT.n0 OUT.t1 180.101
R45 OUT OUT.n0 9.363
R46 B.n0 B.t1 795.301
R47 B.n0 B.t0 216.9
R48 B.n1 B.n0 161.3
R49 B B.n1 0.063
R50 B.n1 B 0.063
R51 a_240_100.t0 a_240_100.t1 60.0005
R52 VN.t4 VN.n1 1914.81
R53 VN.n2 VN.t2 1772.88
R54 VN.n1 VN.t0 1181.48
R55 VN.t2 VN.t4 1059.26
R56 VN.n1 VN.n0 591.4
R57 VN.n2 VN.t3 122.501
R58 VN.n0 VN.t1 122.501
R59 VN VN.n0 38.4338
R60 VN.n3 VN.n2 38.1005
R61 VN VN.n3 0.729667
R62 VN.n3 VN 0.333833
R63 A.n0 A.t1 579.861
R64 A.n0 A.t0 419.195
R65 A.n1 A.n0 161.3
R66 A A.n1 0.063
R67 A.n1 A 0.063
C0 VP OUT 0.23994f
C1 VP nand_0.OUT 0.59969f
C2 VP B 0.07471f
C3 A nand_0.OUT 0.07079f
C4 OUT nand_0.OUT 0.1265f
C5 A B 0.0726f
C6 nand_0.OUT B 0.14344f
C7 VP A 0.12794f
C8 OUT VN 0.36041f
C9 B VN 0.2723f
C10 A VN 0.31571f
C11 VP VN 2.11794f
C12 nand_0.OUT VN 0.57391f
.ends

