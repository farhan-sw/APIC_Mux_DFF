* PEX produced on Sat Apr 12 06:59:30 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from top_level.ext - technology: sky130A

.subckt top_level A B S Clk Q Qi VP VN
X0 mux_0.or_0.nor_0.OUT.t2 mux_0.or_0.B.t2 a_2480_580.t1 VP.t36 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X1 Q.t2 Qi.t3 a_4810_100.t1 VN.t27 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X2 Qi.t0 dff_1.nand_2.B.t3 a_5320_100.t0 VN.t2 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X3 a_2480_580.t0 mux_0.or_0.A.t2 VP.t11 VP.t10 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X4 VP.t3 A.t0 mux_0.and_0.nand_0.OUT.t2 VP.t2 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X5 VP.t9 Qi.t4 Q.t1 VP.t8 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X6 VP.t23 dff_1.nand_2.B.t4 Qi.t1 VP.t22 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X7 mux_0.D.t0 mux_0.or_0.nor_0.OUT.t3 VN.t29 VN.t28 sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X8 dff_1.nand_0.A.t0 mux_0.D.t2 VN.t8 VN.t7 sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X9 mux_0.D.t1 mux_0.or_0.nor_0.OUT.t4 VP.t35 VP.t34 sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X10 dff_1.nand_0.A.t1 mux_0.D.t3 VP.t29 VP.t28 sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X11 mux_0.or_0.B.t1 mux_0.and_0.nand_0.OUT.t3 VN.t19 VN.t18 sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X12 mux_0.or_0.B.t0 mux_0.and_0.nand_0.OUT.t4 VP.t15 VP.t14 sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X13 dff_1.nand_2.B.t1 Clk.t0 a_3790_100.t0 VN.t12 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X14 a_3790_100.t1 dff_1.nand_0.A.t2 VN.t25 VN.t24 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X15 a_4300_100.t0 mux_0.D.t4 VN.t11 VN.t10 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X16 mux_0.and_1.nand_0.OUT.t2 S.t0 a_1550_100.t1 VN.t15 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X17 VP.t31 Clk.t1 dff_1.nand_2.B.t2 VP.t30 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X18 a_1550_100.t0 B.t0 VN.t23 VN.t22 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X19 mux_0.or_0.A.t1 mux_0.and_1.nand_0.OUT.t3 VN.t6 VN.t5 sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X20 dff_1.nand_2.B.t0 dff_1.nand_0.A.t3 VP.t17 VP.t16 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X21 dff_1.nand_3.A.t0 mux_0.D.t5 VP.t13 VP.t12 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X22 VP.t5 S.t1 mux_0.and_1.nand_0.OUT.t1 VP.t4 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X23 mux_0.inverter_0.OUT.t0 S.t2 VN.t14 VN.t13 sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X24 dff_1.nand_3.A.t2 Clk.t2 a_4300_100.t1 VN.t26 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X25 mux_0.and_1.nand_0.OUT.t0 B.t1 VP.t21 VP.t20 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X26 mux_0.or_0.A.t0 mux_0.and_1.nand_0.OUT.t4 VP.t1 VP.t0 sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X27 a_620_100.t0 mux_0.inverter_0.OUT.t2 VN.t1 VN.t0 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X28 a_4810_100.t0 dff_1.nand_3.A.t3 VN.t17 VN.t16 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X29 a_5320_100.t1 Q.t3 VN.t21 VN.t20 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
X30 mux_0.inverter_0.OUT.t1 S.t3 VP.t27 VP.t26 sky130_fd_pr__pfet_01v8 ad=1.35 pd=6.9 as=1.35 ps=6.9 w=3 l=0.15
X31 VP.t19 Clk.t3 dff_1.nand_3.A.t1 VP.t18 sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=0.15
X32 VN.t31 mux_0.or_0.B.t3 mux_0.or_0.nor_0.OUT.t1 VN.t30 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X33 mux_0.and_0.nand_0.OUT.t0 mux_0.inverter_0.OUT.t3 VP.t7 VP.t6 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X34 Qi.t2 Q.t4 VP.t33 VP.t32 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X35 Q.t0 dff_1.nand_3.A.t4 VP.t25 VP.t24 sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.35 ps=6.9 w=3 l=0.15
X36 mux_0.and_0.nand_0.OUT.t1 A.t1 a_620_100.t1 VN.t9 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X37 mux_0.or_0.nor_0.OUT.t0 mux_0.or_0.A.t3 VN.t4 VN.t3 sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.45 ps=2.9 w=1 l=0.15
R0 mux_0.or_0.B.n0 mux_0.or_0.B.t2 586.433
R1 mux_0.or_0.B.n0 mux_0.or_0.B.t3 425.767
R2 mux_0.or_0.B.n1 mux_0.or_0.B.t0 190.534
R3 mux_0.or_0.B.n1 mux_0.or_0.B.t1 180.101
R4 mux_0.or_0.nor_0.B mux_0.or_0.B.n0 161.3
R5 mux_0.or_0.nor_0.B mux_0.or_0.B.n1 32.1755
R6 a_2480_580.t0 a_2480_580.t1 32.8338
R7 mux_0.or_0.nor_0.OUT.n0 mux_0.or_0.nor_0.OUT.t4 660.194
R8 mux_0.or_0.nor_0.OUT.n0 mux_0.or_0.nor_0.OUT.t3 338.861
R9 mux_0.or_0.nor_0.OUT.n2 mux_0.or_0.nor_0.OUT.t2 209.733
R10 mux_0.or_0.nor_0.OUT mux_0.or_0.nor_0.OUT.n0 161.363
R11 mux_0.or_0.nor_0.OUT.n2 mux_0.or_0.nor_0.OUT.n1 156.5
R12 mux_0.or_0.nor_0.OUT.n1 mux_0.or_0.nor_0.OUT.t1 30.0005
R13 mux_0.or_0.nor_0.OUT.n1 mux_0.or_0.nor_0.OUT.t0 30.0005
R14 mux_0.or_0.nor_0.OUT mux_0.or_0.nor_0.OUT.n2 9.363
R15 VP.n54 VP.t34 384.192
R16 VP.t0 VP.n74 384.192
R17 VP.n115 VP.t14 384.192
R18 VP.n20 VP.t8 328.31
R19 VP.t18 VP.n32 328.31
R20 VP.n37 VP.t30 328.31
R21 VP.t28 VP.n49 328.31
R22 VP.t36 VP.n65 328.31
R23 VP.n120 VP.t4 328.31
R24 VP.n104 VP.t2 328.31
R25 VP.n99 VP.t26 328.31
R26 VP.n87 VP.n85 300
R27 VP.n81 VP.n80 300
R28 VP.n103 VP.n79 300
R29 VP.n76 VP.n75 300
R30 VP.n119 VP.n2 300
R31 VP.n67 VP.n66 300
R32 VP.n4 VP.n3 300
R33 VP.n53 VP.n6 300
R34 VP.n8 VP.n7 300
R35 VP.n36 VP.n11 300
R36 VP.n13 VP.n12 300
R37 VP.n19 VP.n15 300
R38 VP.n90 VP.n89 292.5
R39 VP.n95 VP.n94 292.5
R40 VP.n102 VP.n100 292.5
R41 VP.n111 VP.n110 292.5
R42 VP.n118 VP.n116 292.5
R43 VP.n70 VP.n69 292.5
R44 VP.n61 VP.n60 292.5
R45 VP.n52 VP.n50 292.5
R46 VP.n45 VP.n44 292.5
R47 VP.n35 VP.n33 292.5
R48 VP.n28 VP.n27 292.5
R49 VP.n18 VP.n16 292.5
R50 VP.n20 VP.t32 202.575
R51 VP.n32 VP.t24 202.575
R52 VP.n37 VP.t12 202.575
R53 VP.n49 VP.t16 202.575
R54 VP.n54 VP.t28 202.575
R55 VP.n65 VP.t34 202.575
R56 VP.n74 VP.t10 202.575
R57 VP.n120 VP.t0 202.575
R58 VP.t20 VP.n115 202.575
R59 VP.n104 VP.t14 202.575
R60 VP.t6 VP.n99 202.575
R61 VP.n86 VP.t26 202.575
R62 VP.n23 VP.t23 184.375
R63 VP.n82 VP.t3 183.833
R64 VP.n77 VP.t5 183.833
R65 VP.n41 VP.t31 183.833
R66 VP.n9 VP.t19 183.833
R67 VP.n24 VP.t9 183.833
R68 VP.t32 VP.t22 181.619
R69 VP.t8 VP.t24 181.619
R70 VP.t12 VP.t18 181.619
R71 VP.t30 VP.t16 181.619
R72 VP.t10 VP.t36 181.619
R73 VP.t4 VP.t20 181.619
R74 VP.t2 VP.t6 181.619
R75 VP.n98 VP.n97 149.718
R76 VP.n106 VP.n105 149.718
R77 VP.n114 VP.n113 149.718
R78 VP.n122 VP.n121 149.718
R79 VP.n73 VP.n72 149.718
R80 VP.n64 VP.n63 149.718
R81 VP.n56 VP.n55 149.718
R82 VP.n48 VP.n47 149.718
R83 VP.n39 VP.n38 149.718
R84 VP.n31 VP.n30 149.718
R85 VP.n90 VP.n83 149.718
R86 VP.n22 VP.n21 149.718
R87 VP.n89 VP.n88 141.603
R88 VP.n96 VP.n95 140.119
R89 VP.n100 VP.n78 140.119
R90 VP.n112 VP.n111 140.119
R91 VP.n116 VP.n1 140.119
R92 VP.n71 VP.n70 140.119
R93 VP.n62 VP.n61 140.119
R94 VP.n50 VP.n5 140.119
R95 VP.n46 VP.n45 140.119
R96 VP.n33 VP.n10 140.119
R97 VP.n29 VP.n28 140.119
R98 VP.n16 VP.n14 140.119
R99 VP.n88 VP.n87 108.195
R100 VP.n94 VP.n80 98.9005
R101 VP.n103 VP.n102 98.9005
R102 VP.n110 VP.n75 98.9005
R103 VP.n119 VP.n118 98.9005
R104 VP.n69 VP.n66 98.9005
R105 VP.n60 VP.n3 98.9005
R106 VP.n53 VP.n52 98.9005
R107 VP.n44 VP.n7 98.9005
R108 VP.n36 VP.n35 98.9005
R109 VP.n27 VP.n12 98.9005
R110 VP.n19 VP.n18 98.9005
R111 VP.n26 VP.n13 92.5005
R112 VP.n32 VP.n12 92.5005
R113 VP.n34 VP.n11 92.5005
R114 VP.n37 VP.n36 92.5005
R115 VP.n43 VP.n8 92.5005
R116 VP.n49 VP.n7 92.5005
R117 VP.n51 VP.n6 92.5005
R118 VP.n54 VP.n53 92.5005
R119 VP.n59 VP.n4 92.5005
R120 VP.n65 VP.n3 92.5005
R121 VP.n68 VP.n67 92.5005
R122 VP.n74 VP.n66 92.5005
R123 VP.n117 VP.n2 92.5005
R124 VP.n120 VP.n119 92.5005
R125 VP.n109 VP.n76 92.5005
R126 VP.n115 VP.n75 92.5005
R127 VP.n101 VP.n79 92.5005
R128 VP.n104 VP.n103 92.5005
R129 VP.n93 VP.n81 92.5005
R130 VP.n99 VP.n80 92.5005
R131 VP.n85 VP.n84 92.5005
R132 VP.n87 VP.n86 92.5005
R133 VP.n20 VP.n19 92.5005
R134 VP.n17 VP.n15 92.5005
R135 VP.n85 VP.n83 57.2175
R136 VP.n31 VP.n13 57.2175
R137 VP.n38 VP.n11 57.2175
R138 VP.n48 VP.n8 57.2175
R139 VP.n55 VP.n6 57.2175
R140 VP.n64 VP.n4 57.2175
R141 VP.n73 VP.n67 57.2175
R142 VP.n121 VP.n2 57.2175
R143 VP.n114 VP.n76 57.2175
R144 VP.n105 VP.n79 57.2175
R145 VP.n98 VP.n81 57.2175
R146 VP.n21 VP.n15 57.2175
R147 VP.n91 VP.n90 44.5005
R148 VP.n97 VP.n92 44.5005
R149 VP.n107 VP.n106 44.5005
R150 VP.n113 VP.n108 44.5005
R151 VP.n123 VP.n122 44.5005
R152 VP.n72 VP.n0 44.5005
R153 VP.n63 VP.n58 44.5005
R154 VP.n57 VP.n56 44.5005
R155 VP.n47 VP.n42 44.5005
R156 VP.n40 VP.n39 44.5005
R157 VP.n30 VP.n25 44.5005
R158 VP.n23 VP.n22 44.5005
R159 VP.n90 VP.n84 25.6005
R160 VP.n94 VP.n93 19.2005
R161 VP.n102 VP.n101 19.2005
R162 VP.n110 VP.n109 19.2005
R163 VP.n118 VP.n117 19.2005
R164 VP.n69 VP.n68 19.2005
R165 VP.n60 VP.n59 19.2005
R166 VP.n52 VP.n51 19.2005
R167 VP.n44 VP.n43 19.2005
R168 VP.n35 VP.n34 19.2005
R169 VP.n27 VP.n26 19.2005
R170 VP.n18 VP.n17 19.2005
R171 VP.n32 VP.n31 17.6428
R172 VP.n38 VP.n37 17.6428
R173 VP.n49 VP.n48 17.6428
R174 VP.n55 VP.n54 17.6428
R175 VP.n65 VP.n64 17.6428
R176 VP.n74 VP.n73 17.6428
R177 VP.n121 VP.n120 17.6428
R178 VP.n115 VP.n114 17.6428
R179 VP.n105 VP.n104 17.6428
R180 VP.n99 VP.n98 17.6428
R181 VP.n86 VP.n83 17.6428
R182 VP.n21 VP.n20 17.6428
R183 VP.n89 VP.t27 16.4172
R184 VP.n95 VP.t7 16.4172
R185 VP.n100 VP.t15 16.4172
R186 VP.n111 VP.t21 16.4172
R187 VP.n116 VP.t1 16.4172
R188 VP.n70 VP.t11 16.4172
R189 VP.n61 VP.t35 16.4172
R190 VP.n50 VP.t29 16.4172
R191 VP.n45 VP.t17 16.4172
R192 VP.n33 VP.t13 16.4172
R193 VP.n28 VP.t25 16.4172
R194 VP.n16 VP.t33 16.4172
R195 VP.n97 VP.n96 12.2643
R196 VP.n96 VP.n93 12.2643
R197 VP.n106 VP.n78 12.2643
R198 VP.n101 VP.n78 12.2643
R199 VP.n113 VP.n112 12.2643
R200 VP.n112 VP.n109 12.2643
R201 VP.n122 VP.n1 12.2643
R202 VP.n117 VP.n1 12.2643
R203 VP.n72 VP.n71 12.2643
R204 VP.n71 VP.n68 12.2643
R205 VP.n63 VP.n62 12.2643
R206 VP.n62 VP.n59 12.2643
R207 VP.n56 VP.n5 12.2643
R208 VP.n51 VP.n5 12.2643
R209 VP.n47 VP.n46 12.2643
R210 VP.n46 VP.n43 12.2643
R211 VP.n39 VP.n10 12.2643
R212 VP.n34 VP.n10 12.2643
R213 VP.n30 VP.n29 12.2643
R214 VP.n29 VP.n26 12.2643
R215 VP.n22 VP.n14 12.2643
R216 VP.n17 VP.n14 12.2643
R217 VP.n88 VP.n84 9.29594
R218 VP VP.n0 0.729667
R219 VP.n25 VP.n24 0.542167
R220 VP.n40 VP.n9 0.542167
R221 VP.n42 VP.n41 0.542167
R222 VP.n58 VP 0.542167
R223 VP VP.n123 0.542167
R224 VP.n108 VP.n77 0.542167
R225 VP VP.n107 0.542167
R226 VP.n92 VP.n82 0.542167
R227 VP.n57 VP 0.458833
R228 VP VP.n91 0.458833
R229 VP VP.n23 0.333833
R230 VP.n25 VP 0.333833
R231 VP VP.n40 0.333833
R232 VP.n42 VP 0.333833
R233 VP VP.n57 0.333833
R234 VP.n58 VP 0.333833
R235 VP VP.n0 0.333833
R236 VP.n123 VP 0.333833
R237 VP.n108 VP 0.333833
R238 VP.n107 VP 0.333833
R239 VP.n92 VP 0.333833
R240 VP.n91 VP 0.333833
R241 VP.n24 VP 0.188
R242 VP VP.n9 0.188
R243 VP.n41 VP 0.188
R244 VP.n77 VP 0.188
R245 VP.n82 VP 0.188
R246 Qi.n0 Qi.t4 795.301
R247 Qi.n0 Qi.t3 216.9
R248 Qi.n3 Qi.t0 196.101
R249 Qi.n3 Qi.n2 183.718
R250 Qi.n1 Qi.n0 161.3
R251 Qi.n4 Qi.n1 21.688
R252 Qi.n2 Qi.t1 16.4172
R253 Qi.n2 Qi.t2 16.4172
R254 Qi.n4 Qi.n3 9.3005
R255 Qi Qi.n4 0.188
R256 Qi.n1 Qi 0.063
R257 a_4810_100.t0 a_4810_100.t1 60.0005
R258 Q.n2 Q.t4 579.861
R259 Q.n2 Q.t3 419.195
R260 Q.n1 Q.t2 196.101
R261 Q.n1 Q.n0 183.718
R262 Q.n3 Q.n2 161.3
R263 Q.n0 Q.t1 16.4172
R264 Q.n0 Q.t0 16.4172
R265 Q.n3 Q 10.0943
R266 Q Q.n1 9.363
R267 Q.n3 Q 0.59425
R268 Q Q.n3 0.063
R269 VN.n12 VN.t28 2240.74
R270 VN.t5 VN.n20 2240.74
R271 VN.n31 VN.t18 2240.74
R272 VN.n1 VN.t27 1914.81
R273 VN.t26 VN.n5 1914.81
R274 VN.n6 VN.t12 1914.81
R275 VN.t7 VN.n11 1914.81
R276 VN.t30 VN.n18 1914.81
R277 VN.n32 VN.t15 1914.81
R278 VN.n26 VN.t9 1914.81
R279 VN.n25 VN.t13 1914.81
R280 VN.n21 VN.t13 1772.88
R281 VN.n1 VN.t20 1181.48
R282 VN.n5 VN.t16 1181.48
R283 VN.n6 VN.t10 1181.48
R284 VN.n11 VN.t24 1181.48
R285 VN.n12 VN.t7 1181.48
R286 VN.n18 VN.t28 1181.48
R287 VN.n20 VN.t3 1181.48
R288 VN.n32 VN.t5 1181.48
R289 VN.t22 VN.n31 1181.48
R290 VN.n26 VN.t18 1181.48
R291 VN.t0 VN.n25 1181.48
R292 VN.t20 VN.t2 1059.26
R293 VN.t27 VN.t16 1059.26
R294 VN.t10 VN.t26 1059.26
R295 VN.t12 VN.t24 1059.26
R296 VN.t3 VN.t30 1059.26
R297 VN.t15 VN.t22 1059.26
R298 VN.t9 VN.t0 1059.26
R299 VN.n25 VN.n24 591.4
R300 VN.n27 VN.n26 591.4
R301 VN.n31 VN.n30 591.4
R302 VN.n33 VN.n32 591.4
R303 VN.n20 VN.n19 591.4
R304 VN.n18 VN.n17 591.4
R305 VN.n13 VN.n12 591.4
R306 VN.n11 VN.n10 591.4
R307 VN.n7 VN.n6 591.4
R308 VN.n5 VN.n4 591.4
R309 VN.n2 VN.n1 591.4
R310 VN.n15 VN.t31 173.4
R311 VN.n21 VN.t14 122.501
R312 VN.n24 VN.t1 122.501
R313 VN.n27 VN.t19 122.501
R314 VN.n30 VN.t23 122.501
R315 VN.n33 VN.t6 122.501
R316 VN.n19 VN.t4 122.501
R317 VN.n17 VN.t29 122.501
R318 VN.n13 VN.t8 122.501
R319 VN.n10 VN.t25 122.501
R320 VN.n7 VN.t11 122.501
R321 VN.n4 VN.t17 122.501
R322 VN.n2 VN.t21 122.501
R323 VN VN.n2 38.4338
R324 VN.n22 VN.n21 38.1005
R325 VN.n24 VN.n23 38.1005
R326 VN.n28 VN.n27 38.1005
R327 VN.n30 VN.n29 38.1005
R328 VN.n34 VN.n33 38.1005
R329 VN.n19 VN.n0 38.1005
R330 VN.n17 VN.n16 38.1005
R331 VN.n14 VN.n13 38.1005
R332 VN.n10 VN.n9 38.1005
R333 VN.n8 VN.n7 38.1005
R334 VN.n4 VN.n3 38.1005
R335 VN.n3 VN 0.729667
R336 VN.n8 VN 0.729667
R337 VN.n9 VN 0.729667
R338 VN.n29 VN 0.729667
R339 VN.n23 VN 0.729667
R340 VN.n16 VN 0.542167
R341 VN.n15 VN.n0 0.542167
R342 VN VN.n34 0.542167
R343 VN VN.n28 0.542167
R344 VN.n14 VN 0.458833
R345 VN VN.n22 0.458833
R346 VN.n3 VN 0.333833
R347 VN VN.n8 0.333833
R348 VN.n9 VN 0.333833
R349 VN VN.n14 0.333833
R350 VN.n16 VN 0.333833
R351 VN VN.n0 0.333833
R352 VN.n34 VN 0.333833
R353 VN.n29 VN 0.333833
R354 VN.n28 VN 0.333833
R355 VN.n23 VN 0.333833
R356 VN.n22 VN 0.333833
R357 VN VN.n15 0.188
R358 dff_1.nand_2.B.n0 dff_1.nand_2.B.t4 795.301
R359 dff_1.nand_2.B.n0 dff_1.nand_2.B.t3 216.9
R360 dff_1.nand_2.B.n2 dff_1.nand_2.B.t1 196.101
R361 dff_1.nand_2.B.n2 dff_1.nand_2.B.n1 183.718
R362 dff_1.nand_2.B dff_1.nand_2.B.n0 161.3
R363 dff_1.nand_2.B dff_1.nand_2.B.n2 32.5505
R364 dff_1.nand_2.B.n1 dff_1.nand_2.B.t2 16.4172
R365 dff_1.nand_2.B.n1 dff_1.nand_2.B.t0 16.4172
R366 a_5320_100.t0 a_5320_100.t1 60.0005
R367 mux_0.or_0.A.n0 mux_0.or_0.A.t2 579.861
R368 mux_0.or_0.A.n0 mux_0.or_0.A.t3 419.195
R369 mux_0.or_0.A.n1 mux_0.or_0.A.t0 190.534
R370 mux_0.or_0.A.n1 mux_0.or_0.A.t1 180.101
R371 mux_0.or_0.nor_0.A mux_0.or_0.A.n0 161.363
R372 mux_0.and_1.inverter_0.OUT mux_0.or_0.A.n1 9.35606
R373 mux_0.and_1.inverter_0.OUT mux_0.or_0.nor_0.A 0.6255
R374 A.n0 A.t0 795.301
R375 A.n0 A.t1 216.9
R376 A A.n0 161.363
R377 mux_0.and_0.nand_0.OUT.n0 mux_0.and_0.nand_0.OUT.t4 660.194
R378 mux_0.and_0.nand_0.OUT.n0 mux_0.and_0.nand_0.OUT.t3 338.861
R379 mux_0.and_0.nand_0.OUT.n2 mux_0.and_0.nand_0.OUT.t1 196.101
R380 mux_0.and_0.nand_0.OUT.n2 mux_0.and_0.nand_0.OUT.n1 183.718
R381 mux_0.and_0.nand_0.OUT mux_0.and_0.nand_0.OUT.n0 161.3
R382 mux_0.and_0.nand_0.OUT.n1 mux_0.and_0.nand_0.OUT.t2 16.4172
R383 mux_0.and_0.nand_0.OUT.n1 mux_0.and_0.nand_0.OUT.t0 16.4172
R384 mux_0.and_0.nand_0.OUT mux_0.and_0.nand_0.OUT.n2 9.363
R385 mux_0.D.n1 mux_0.D.t3 660.194
R386 mux_0.D.n0 mux_0.D.t5 579.861
R387 mux_0.D.n0 mux_0.D.t4 419.195
R388 mux_0.D.n1 mux_0.D.t2 338.861
R389 mux_0.D.n2 mux_0.D.t1 190.534
R390 mux_0.D.n2 mux_0.D.t0 180.101
R391 dff_1.inverter_1.A mux_0.D.n1 161.3
R392 dff_1.nand_1.A mux_0.D.n0 161.3
R393 dff_1.inverter_1.A dff_1.nand_1.A 21.3755
R394 mux_0.or_0.inverter_0.OUT mux_0.D.n2 9.363
R395 mux_0.or_0.inverter_0.OUT dff_1.inverter_1.A 0.688
R396 dff_1.nand_0.A.n0 dff_1.nand_0.A.t3 579.861
R397 dff_1.nand_0.A.n0 dff_1.nand_0.A.t2 419.195
R398 dff_1.nand_0.A.n1 dff_1.nand_0.A.t1 190.534
R399 dff_1.nand_0.A.n1 dff_1.nand_0.A.t0 180.101
R400 dff_1.nand_0.A dff_1.nand_0.A.n0 161.363
R401 dff_1.nand_0.A dff_1.nand_0.A.n1 9.35606
R402 Clk.n1 Clk.t1 795.301
R403 Clk.n0 Clk.t3 795.301
R404 Clk.n1 Clk.t0 216.9
R405 Clk.n0 Clk.t2 216.9
R406 Clk Clk.n0 161.363
R407 Clk.n2 Clk.n1 161.3
R408 Clk.n3 Clk 20.0005
R409 Clk.n3 Clk 1.90675
R410 Clk.n2 Clk 1.40675
R411 Clk Clk.n2 0.063
R412 Clk Clk.n3 0.063
R413 a_3790_100.t0 a_3790_100.t1 60.0005
R414 a_4300_100.t0 a_4300_100.t1 60.0005
R415 S.n0 S.t1 795.301
R416 S.n2 S.t3 660.194
R417 S.n2 S.t2 338.861
R418 S.n0 S.t0 216.9
R419 S.n3 S.n2 161.3
R420 S.n1 S.n0 161.3
R421 S.n3 S.n1 23.7817
R422 S.n1 S 0.063
R423 S S.n3 0.063
R424 a_1550_100.t0 a_1550_100.t1 60.0005
R425 mux_0.and_1.nand_0.OUT.n0 mux_0.and_1.nand_0.OUT.t4 660.194
R426 mux_0.and_1.nand_0.OUT.n0 mux_0.and_1.nand_0.OUT.t3 338.861
R427 mux_0.and_1.nand_0.OUT.n2 mux_0.and_1.nand_0.OUT.t2 196.101
R428 mux_0.and_1.nand_0.OUT.n2 mux_0.and_1.nand_0.OUT.n1 183.718
R429 mux_0.and_1.nand_0.OUT mux_0.and_1.nand_0.OUT.n0 161.3
R430 mux_0.and_1.nand_0.OUT.n1 mux_0.and_1.nand_0.OUT.t1 16.4172
R431 mux_0.and_1.nand_0.OUT.n1 mux_0.and_1.nand_0.OUT.t0 16.4172
R432 mux_0.and_1.nand_0.OUT mux_0.and_1.nand_0.OUT.n2 9.363
R433 B.n0 B.t1 579.861
R434 B.n0 B.t0 419.195
R435 B.n1 B.n0 161.3
R436 B B.n1 13.9693
R437 B.n1 B 0.063
R438 dff_1.nand_3.A.n0 dff_1.nand_3.A.t4 579.861
R439 dff_1.nand_3.A.n0 dff_1.nand_3.A.t3 419.195
R440 dff_1.nand_3.A.n2 dff_1.nand_3.A.t2 196.101
R441 dff_1.nand_3.A.n2 dff_1.nand_3.A.n1 183.718
R442 dff_1.nand_3.A dff_1.nand_3.A.n0 161.3
R443 dff_1.nand_3.A.n1 dff_1.nand_3.A.t1 16.4172
R444 dff_1.nand_3.A.n1 dff_1.nand_3.A.t0 16.4172
R445 dff_1.nand_3.A dff_1.nand_3.A.n2 9.363
R446 mux_0.inverter_0.OUT.n0 mux_0.inverter_0.OUT.t3 579.861
R447 mux_0.inverter_0.OUT.n0 mux_0.inverter_0.OUT.t2 419.195
R448 mux_0.inverter_0.OUT.n1 mux_0.inverter_0.OUT.t1 190.534
R449 mux_0.inverter_0.OUT.n1 mux_0.inverter_0.OUT.t0 180.101
R450 mux_0.inverter_0.OUT mux_0.inverter_0.OUT.n0 161.363
R451 mux_0.inverter_0.OUT mux_0.inverter_0.OUT.n1 9.35606
R452 a_620_100.t0 a_620_100.t1 60.0005
C0 dff_1.nand_0.A VP 0.48118f
C1 mux_0.and_1.nand_0.OUT B 0.08079f
C2 mux_0.and_0.nand_0.OUT A 0.14419f
C3 Q dff_1.nand_3.A 0.08239f
C4 dff_1.nand_2.B Qi 0.61525f
C5 VP Qi 0.51323f
C6 mux_0.and_0.nand_0.OUT S 0.03678f
C7 B Clk 0.01528f
C8 mux_0.inverter_0.OUT VP 0.49374f
C9 mux_0.inverter_0.OUT B 0.03505f
C10 VP A 0.07132f
C11 S VP 0.19299f
C12 B A 0.35798f
C13 S B 0.66535f
C14 dff_1.nand_3.A Clk 0.14797f
C15 Q Qi 0.43472f
C16 dff_1.nand_3.A Qi 0.08746f
C17 mux_0.and_0.nand_0.OUT VP 0.56285f
C18 mux_0.or_0.nor_0.OUT Clk 0.12816f
C19 mux_0.and_1.nand_0.OUT Clk 0.05619f
C20 mux_0.and_0.nand_0.OUT B 0.13823f
C21 dff_1.nand_0.A Clk 0.25414f
C22 VP dff_1.nand_2.B 0.51872f
C23 mux_0.inverter_0.OUT Clk 0.1155f
C24 VP B 0.1252f
C25 mux_0.and_1.nand_0.OUT S 0.17378f
C26 A Clk 0.03473f
C27 S Clk 0.05049f
C28 mux_0.inverter_0.OUT A 0.23022f
C29 Q dff_1.nand_2.B 0.22377f
C30 VP Q 0.78744f
C31 mux_0.inverter_0.OUT S 0.17868f
C32 dff_1.nand_3.A dff_1.nand_2.B 0.12032f
C33 VP dff_1.nand_3.A 0.62333f
C34 S A 0.13813f
C35 mux_0.and_0.nand_0.OUT Clk 0.12121f
C36 VP mux_0.or_0.nor_0.OUT 0.29377f
C37 mux_0.and_1.nand_0.OUT VP 0.54338f
C38 mux_0.inverter_0.OUT mux_0.and_0.nand_0.OUT 0.08389f
C39 dff_1.nand_2.B Clk 0.45049f
C40 dff_1.nand_0.A dff_1.nand_2.B 0.08985f
C41 VP Clk 1.39606f
C42 Q VN 0.5023f
C43 Qi VN 1.01243f
C44 Clk VN 0.86642f
C45 B VN 0.61957f
C46 A VN 0.29322f
C47 S VN 1.68603f
C48 VP VN 12.5509f
C49 dff_1.nand_2.B VN 0.99398f
C50 dff_1.nand_3.A VN 0.43673f
C51 dff_1.nand_0.A VN 0.49658f
C52 mux_0.or_0.nor_0.OUT VN 0.68172f
C53 mux_0.and_1.nand_0.OUT VN 0.53204f
C54 mux_0.and_0.nand_0.OUT VN 0.46924f
C55 mux_0.inverter_0.OUT VN 0.50204f
.ends

