magic
tech sky130A
magscale 1 2
timestamp 1744431535
<< nwell >>
rect 3130 540 3170 1220
<< metal1 >>
rect 0 1220 30 1280
rect 3130 1220 3170 1280
rect 30 750 3250 760
rect 30 720 3180 750
rect 3170 690 3180 720
rect 3240 690 3250 750
rect 3170 680 3250 690
rect 5210 660 5290 670
rect 5210 600 5220 660
rect 5280 650 5290 660
rect 5460 660 5540 670
rect 5460 650 5470 660
rect 5280 610 5470 650
rect 5280 600 5290 610
rect 5210 590 5290 600
rect 5460 600 5470 610
rect 5530 650 5540 660
rect 5530 610 5560 650
rect 5530 600 5540 610
rect 5460 590 5540 600
rect 5210 520 5290 530
rect 5210 460 5220 520
rect 5280 460 5290 520
rect 30 420 70 460
rect 3100 420 3170 460
rect 5210 450 5290 460
rect 5460 520 5540 530
rect 5460 460 5470 520
rect 5530 510 5540 520
rect 5530 470 5560 510
rect 5530 460 5540 470
rect 5460 450 5540 460
rect 30 320 70 360
rect 3170 350 3250 360
rect 3170 290 3180 350
rect 3240 290 3250 350
rect 3170 280 3250 290
rect 30 240 70 280
rect 0 0 30 60
rect 3130 0 3170 60
<< via1 >>
rect 3180 690 3240 750
rect 5220 600 5280 660
rect 5470 600 5530 660
rect 5220 460 5280 520
rect 5470 460 5530 520
rect 3180 290 3240 350
<< metal2 >>
rect 3170 750 3250 760
rect 3170 690 3180 750
rect 3240 690 3250 750
rect 3170 680 3250 690
rect 3190 360 3230 680
rect 5210 660 5290 670
rect 5210 600 5220 660
rect 5280 600 5290 660
rect 5210 590 5290 600
rect 5460 660 5540 670
rect 5460 600 5470 660
rect 5530 600 5540 660
rect 5460 590 5540 600
rect 5230 530 5270 590
rect 5210 520 5290 530
rect 5210 460 5220 520
rect 5280 460 5290 520
rect 5210 450 5290 460
rect 5460 520 5540 530
rect 5460 460 5470 520
rect 5530 460 5540 520
rect 5460 450 5540 460
rect 3170 350 3250 360
rect 3170 290 3180 350
rect 3240 290 3250 350
rect 3170 280 3250 290
use dff  dff_1
timestamp 1744388325
transform 1 0 3170 0 1 0
box 0 0 2420 1280
use mux  mux_0
timestamp 1744416606
transform 1 0 0 0 1 0
box 0 0 3171 1280
<< labels >>
flabel metal1 30 420 30 460 1 FreeSans 560 0 0 0 S
port 3 n
flabel metal1 30 320 30 360 1 FreeSans 560 0 0 0 A
port 1 n
flabel metal1 30 240 30 280 1 FreeSans 560 0 0 0 B
port 2 n
flabel metal1 30 720 30 760 1 FreeSans 560 0 0 0 Clk
port 4 n
flabel metal1 5560 610 5560 650 1 FreeSans 560 0 0 0 Q
port 5 n
flabel metal1 5560 470 5560 510 1 FreeSans 560 0 0 0 Qi
port 6 n
flabel metal1 0 1220 0 1280 3 FreeSans 560 0 0 0 VP
port 7 e
flabel metal1 0 0 0 60 3 FreeSans 560 0 0 0 VN
port 8 e
<< end >>
