magic
tech sky130A
timestamp 1744374832
<< nwell >>
rect -105 220 150 560
<< nmos >>
rect 0 0 15 100
rect 65 0 80 100
<< pmos >>
rect 0 240 15 540
rect 65 240 80 540
<< ndiff >>
rect -45 85 0 100
rect -45 15 -35 85
rect -15 15 0 85
rect -45 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
<< pdiff >>
rect -45 525 0 540
rect -45 455 -35 525
rect -15 455 0 525
rect -45 425 0 455
rect -45 355 -35 425
rect -15 355 0 425
rect -45 325 0 355
rect -45 255 -35 325
rect -15 255 0 325
rect -45 240 0 255
rect 15 525 65 540
rect 15 455 30 525
rect 50 455 65 525
rect 15 425 65 455
rect 15 355 30 425
rect 50 355 65 425
rect 15 325 65 355
rect 15 255 30 325
rect 50 255 65 325
rect 15 240 65 255
rect 80 525 130 540
rect 80 455 95 525
rect 115 455 130 525
rect 80 425 130 455
rect 80 355 95 425
rect 115 355 130 425
rect 80 325 130 355
rect 80 255 95 325
rect 115 255 130 325
rect 80 240 130 255
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
rect 95 15 115 85
<< pdiffc >>
rect -35 455 -15 525
rect -35 355 -15 425
rect -35 255 -15 325
rect 30 455 50 525
rect 30 355 50 425
rect 30 255 50 325
rect 95 455 115 525
rect 95 355 115 425
rect 95 255 115 325
<< psubdiff >>
rect -85 85 -45 100
rect -85 15 -75 85
rect -55 15 -45 85
rect -85 0 -45 15
<< nsubdiff >>
rect -85 525 -45 540
rect -85 455 -75 525
rect -55 455 -45 525
rect -85 425 -45 455
rect -85 355 -75 425
rect -55 355 -45 425
rect -85 325 -45 355
rect -85 255 -75 325
rect -55 255 -45 325
rect -85 240 -45 255
<< psubdiffcont >>
rect -75 15 -55 85
<< nsubdiffcont >>
rect -75 455 -55 525
rect -75 355 -55 425
rect -75 255 -55 325
<< poly >>
rect 0 540 15 555
rect 65 540 80 555
rect 0 215 15 240
rect 65 215 80 240
rect -40 205 15 215
rect -40 185 -30 205
rect -10 185 15 205
rect -40 175 15 185
rect 40 205 80 215
rect 40 185 50 205
rect 70 185 80 205
rect 40 175 80 185
rect 0 100 15 175
rect 65 100 80 175
rect 0 -15 15 0
rect 65 -15 80 0
<< polycont >>
rect -30 185 -10 205
rect 50 185 70 205
<< locali >>
rect -35 585 -15 590
rect -35 530 -15 565
rect -85 525 -5 530
rect -85 455 -75 525
rect -55 455 -35 525
rect -15 455 -5 525
rect -85 450 -5 455
rect 20 525 60 530
rect 20 455 30 525
rect 50 455 60 525
rect 20 450 60 455
rect 85 525 125 530
rect 85 455 95 525
rect 115 455 125 525
rect 85 450 125 455
rect -35 430 -15 450
rect 30 430 50 450
rect 95 430 115 450
rect -85 425 -5 430
rect -85 355 -75 425
rect -55 355 -35 425
rect -15 355 -5 425
rect -85 350 -5 355
rect 20 425 60 430
rect 20 355 30 425
rect 50 355 60 425
rect 20 350 60 355
rect 85 425 125 430
rect 85 355 95 425
rect 115 355 125 425
rect 85 350 125 355
rect -35 330 -15 350
rect 30 330 50 350
rect 95 330 115 350
rect -85 325 -5 330
rect -85 255 -75 325
rect -55 255 -35 325
rect -15 255 -5 325
rect -85 250 -5 255
rect 20 325 60 330
rect 20 255 30 325
rect 50 255 60 325
rect 20 250 60 255
rect 85 325 125 330
rect 85 255 95 325
rect 115 255 125 325
rect 85 250 125 255
rect -40 205 0 215
rect -40 185 -30 205
rect -10 185 0 205
rect -40 175 0 185
rect 40 205 80 215
rect 40 185 50 205
rect 70 185 80 205
rect 40 175 80 185
rect 105 155 125 250
rect 85 145 125 155
rect 85 135 95 145
rect 30 125 95 135
rect 115 125 125 145
rect 30 115 125 125
rect 30 90 50 115
rect -85 85 -5 90
rect -85 15 -75 85
rect -55 15 -35 85
rect -15 15 -5 85
rect -85 10 -5 15
rect 20 85 60 90
rect 20 15 30 85
rect 50 15 60 85
rect 20 10 60 15
rect 85 85 125 90
rect 85 15 95 85
rect 115 15 125 85
rect 85 10 125 15
rect -35 -25 -15 10
rect 95 -25 115 10
<< viali >>
rect -35 565 -15 585
rect -30 185 -10 205
rect 50 185 70 205
rect 95 125 115 145
rect -35 -45 -15 -25
rect 95 -45 115 -25
<< metal1 >>
rect -105 585 150 590
rect -105 565 -35 585
rect -15 565 150 585
rect -105 560 150 565
rect -40 205 0 215
rect -40 185 -30 205
rect -10 185 0 205
rect -40 175 0 185
rect 40 205 80 215
rect 40 185 50 205
rect 70 185 80 205
rect 40 175 80 185
rect 85 145 125 155
rect 85 125 95 145
rect 115 125 125 145
rect 85 115 125 125
rect -105 -25 150 -20
rect -105 -45 -35 -25
rect -15 -45 95 -25
rect 115 -45 150 -25
rect -105 -50 150 -45
<< labels >>
flabel metal1 -40 175 -40 215 1 FreeSans 200 0 0 0 A
port 1 n
flabel metal1 -105 560 -105 590 3 FreeSans 200 0 0 0 VP
port 4 e
flabel metal1 -105 -50 -105 -20 3 FreeSans 200 0 0 0 VN
port 5 e
flabel metal1 40 175 40 215 1 FreeSans 200 0 0 0 B
port 2 n
flabel metal1 125 115 125 155 1 FreeSans 200 0 0 0 OUT
port 3 n
<< end >>
